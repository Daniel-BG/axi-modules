package am_data_types is
    type am_last_policy_t is (PASS_ZERO, PASS_ONE, OR_ALL, AND_ALL); 
end package;

package body am_data_types is

end am_data_types;